////////////////////////////////////////////////////////////////////////
// Developer Name : Mohsan Naeem 
// Contact info   : mohsannaeem1576@gmail.com
// Module Name    : dummy_seq_pkg
// Description    : Dummy seq_pkg which can be used to create new seq_pkg
///////////////////////////////////////////////////////////////////////
package dummy_seq_pkg;
	import uvm_pkg::*;
	`include "uvm_macros.svh"
	`include "dummy_seq_item.sv"
	`include "dummy_base_sequence.sv"
endpackage