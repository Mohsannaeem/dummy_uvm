////////////////////////////////////////////////////////////////////////
// Developer Name : Mohsan Naeem 
// Contact info   : mohsannaeem1576@gmail.com
// Module Name    : dummy_test_pkg
// Description    : Dummy Test Package which can be used to create new test pkg
///////////////////////////////////////////////////////////////////////
package dummy_test_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    import dummy_seq_pkg::*;
    import dummy_env_pkg::*;
    `include "dummy_base_test.sv"
endpackage